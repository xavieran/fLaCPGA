module RiceFeeder(input iClock,
						input iReset,
						input iEnable,
						input iData,
						output signed [31:0] oData);
						

reg state;






endmodule
