/* The optimal rice parameter can be estimated from the expectation of the sequence
   of numbers as log(|E|, 2) according to  Weinberger (1996)
   */


module CalculateOptimalRice (

    );



endmodule